
`timescale 1ns / 1ps

module tb_fpga;
    integer         error_count = 0;

	reg 			rst_n_0;
	reg 			rst_n_1;

	reg 			D_0	;
	reg 			S_0	;	
	reg 			D_1	;
	reg 			S_1	;	

//#################################################################################################	
//FPGA
//#################################################################################################		
	
//#################################################################################################	
//BFM IEEE1355
//#################################################################################################	
	bfm_ieee1355	
	#(
		.G_MAX_BIT_RATE_Mbs	(100)
	)	
	bfm_ieee1355_0
	(  
		.rst_n				( rst_n_0 ),

		.D_in				( D_0 ),
		.S_in				( S_0 ),
		
		.D_out				( D_1 ),
		.S_out				( S_1 )
    );	

	bfm_ieee1355	
	#(
		.G_MAX_BIT_RATE_Mbs	(100)
	)	
	bfm_ieee1355_1
	(  
		.rst_n				( rst_n_1 ),

		.D_in				( D_1 ),
		.S_in				( S_1 ),
		
		.D_out				( D_0 ),
		.S_out				( S_0 )
    );	
	
	
//#################################################################################################	
//
//#################################################################################################		
   initial
      $timeformat (-9, 3, " ns", 13);	

	initial
	begin
		#0  	rst_n_0 = 1'b0;
		#0  	rst_n_1 = 1'b0;

		#705    rst_n_0 = 1'b1;	
		#151 	rst_n_1 = 1'b1;				
	end




	  

//#################################################################################################	
//TEST SCRIPT
//#################################################################################################	
	initial
	begin
		$display("TEST STARTED");
		
		#50000;

		bfm_ieee1355_0.insert_10b( 10'b1111000011);		
		#50000;
		
		bfm_ieee1355_0.insert_10b( 10'b0011001100);
		bfm_ieee1355_0.insert_10b( 10'b1111111111);
		bfm_ieee1355_0.insert_10b( 10'b0000000000);		
		bfm_ieee1355_0.insert_10b( 10'b1111111111);
		bfm_ieee1355_0.insert_10b( 10'b0000000000);
		bfm_ieee1355_0.insert_10b( 10'b1111111111);
		
		bfm_ieee1355_1.fifo_rx.wait_fill_level(6);	
		#50000;		
		
		
		
		if ( error_count==0 ) $display("TEST PASSED");
		else                  $display("TEST FAILED : %d ERRORS", error_count );
		
		$finish;
	end

endmodule

